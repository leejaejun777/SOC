module weight()

endmodule
